
interface adder_if (clk);
input bit clk ;
logic [3:0] a,b ;
logic [4:0] c ;
 adder_top
endinterface : adder_if // Interface